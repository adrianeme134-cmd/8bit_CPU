`timescale 1ns / 1ps


module CPU_Core(
    input wire clk,
    input wire rst,
    output wire [7:0] ALU_Data,
    output wire [5:0] Current_state,
    output wire [7:0] PC,
    output wire [7:0] REG1,
    output wire [7:0] REG2,
    output wire [15:0] Current_fetch,
    output wire IRWrite_Top,
    output wire MemWrite_Top,
    output wire MemRead_Top,
    output wire PC_en_Top,
    output wire RegWrite_Top

    
    );
    
    // Define instruction opcodes
    parameter addi = 4'b0000;
    parameter add = 4'b0001;
    parameter lw = 4'b0010;
    parameter subi = 4'b0011;
    parameter sub = 4'b0100;
    parameter beq  = 4'b0101;
    parameter bne  = 4'b0110;
    parameter slt = 4'b0111;
    parameter slti = 4'b1000;
    parameter jump = 4'b1001;
    parameter sw = 4'b1010;
    parameter sra = 4'b1011;
    parameter sll = 4'b1100;
    parameter HLT = 4'b1101;
    parameter bitNAND = 4'b1110;
    parameter blt = 4'b1111;
    
     
    // Decoder Interface
    wire [2:0] Register_Destination;// wire that connects to Register file
    wire [2:0] Register_1_operand; // wire that connects to Register file
    wire [2:0] Register_2_operand; // wire that connects to Register file
    wire ALUsrc; //Flag, 1 for immediate instructions 0 for Reg to reg instructions
    wire [3:0] instr_Opcode; //Opcode generated from instruction
    wire [15:0] Fetch; // coming from IR
    wire [5:0] immediate; // acutal immediate value
    wire Is_immediate; // use immediate field
    wire signed_immediate; // will sign extend if immediate needs to be signed or leave as is if unsigned
    wire [11:0] jmp_addr; // We can jump up to 4KB
    wire [3:0] ALUOp; // 4 bit ALU wire Operation code coming out to ALU
    

    
    //Immediate Extension for signed/unsigned
    wire [7:0] extended_immediate;
    
    //sign extenstion unit will choose between unsigned and signed int and will zero extend for unsigned and sign extend for signed
    assign extended_immediate = (signed_immediate) ? {{2{immediate[5]}},immediate} : {{2{1'b0}},immediate};
    
    //ALU Interface
    wire [7:0] ALU_Out_Sequential;
    wire overflow;
    wire less_than_flag;
    wire is_equal;
    wire zero_flag;
    wire [7:0] HI;
    wire [7:0] LO;
    wire [7:0] B;
    wire [7:0] A;
    
    
    // Program counter interface
    wire [7:0] pc; // register that comes out of program counter module
    wire [7:0] next_pc_value; //Branching and jumping target PC (target Address)
  
    
    (* keep_hierarchy = "yes" *)
    Decoder Decoder_module(
    .Fetch(Fetch), // Driven by IR DONE
    .Register_Destination(Register_Destination), // Outputting reg destination DONE
    .Register_1_operand(Register_1_operand), // Outputting Reg 1 operand DONE
    .Register_2_operand(Register_2_operand), // Outputting Reg 2 operand DONE
    .instr_Opcode(instr_Opcode), // Outputting 4 bit instruction Opcode DONE
    .Is_immediate(Is_immediate), // outputting immediate flag for sign extension if needed DONE
    .immediate(immediate), // outputting 6 bit immediate value DONE
    .ALUOp(ALUOp), // Outputting 4 bit ALU op signal DONE
    .jmp_addr(jmp_addr), // outputting 12 bit address field for jump instr DONE
    .signed_immediate(signed_immediate) // outputting if it is a signed or unsigned immediate DONE
    );
    
    
    // FSM Interface 
    wire MemWrite; // Control flag to write to RAM
    wire MemRead; // Flag to read from RAM
    wire IRWrite; //Flag to write to Instruction Register
    wire PC_en; // Signal coming in from FSM to enable PC
    wire RegWrite; // Signal generated by FSM to be used by Register file
    wire ALU_Enable;
    wire [5:0] State; // Probing FSM state register in top level
    
    //PC Interfrace
    reg branch_en; // Signal for FSM 
   
    
    // Datapath mux that decides branching/logic
    always @(*) begin
        branch_en = 1'b0;
        case(instr_Opcode)
            beq: branch_en = (is_equal) ? 1'b1 : 1'b0;
            bne: branch_en = (~is_equal) ? 1'b1 : 1'b0;
            jump: branch_en = 1'b1;
            blt: branch_en = (less_than_flag) ? 1'b1 : 1'b0;
        endcase  
    end
    
    (* keep_hierarchy = "yes" *)
    FSM Control_Logic_Module(
    .clk(clk), // Global clock DONE
    .rst(rst), // Global rst DONE
    .Opcode(instr_Opcode), // instruction opcode driven by decoder DONE
    .MemWrite(MemWrite), // Outputting Write signal to RAM DONE
    .RegWrite(RegWrite), // Outputting RegWrite signal DONE
    .MemRead(MemRead), // Outputting MemRead signal DONE
    .PCWrite(PC_en), // Outputting PC_en signal DONE
    .IRWrite(IRWrite), // Outputting IRWrite signal DONE
    .ALU_Enable(ALU_Enable),
    .State(State) // Probing state for top level module
    );
    
        
    
   // IR interface 
   (* keep_hierarchy = "yes" *) 
   Instruction_Register IR(
   .clk(clk), // Global clock DONE
   .IR_Write(IRWrite), // IR_Write will be driven by FSM DONE
   .pc_add(pc), // addr will be driven by PC DONE
   .Fetch(Fetch) // will output the 16 bit instruction DONE
   );


    // Program counter will start at byte 0 and increment each clk when FSM asserts signal
    (* keep_hierarchy = "yes" *)
    PC program_counter_module(
    .clk(clk), // Global clock DONE
    .rst(rst), // Global rst DONE
    .PC_en(PC_en), // FSM generated driven signal DONE
    .jump_en(branch_en), // this signal has to come from datapath MUX DONE
    .next_pc_value(extended_immediate), // comes from decoder as unsigned immediate DONE
    .pc(pc) // current addr value DONE
    );


    // assign Fetch = {instruction_byte[pc+1],instruction_byte[pc]}; this is a mistake and we cannot do this because program counter signals are not stable and will flick through states
    // Fetch must be a reg implying it must be clocked for signal stability

   
   // Register file Interface
    wire [7:0] register_1_data; // Outputting Reg 1 data from Register file at all times (combinational read)
    wire [7:0] register_2_data; // Outputting Reg 2 data from Register file at all times (combinational read)
    wire [7:0] data_in_REG; // Wire from data driven by RAM or ALU
    wire [7:0] RAM_data_out;
    
    assign data_in_REG = (instr_Opcode == lw) ? RAM_data_out : ALU_Out_Sequential; // chooses between RAM or ALU as data going in
    
    
    (* keep_hierarchy = "yes" *)
    Register_file Reg_module(
    .rst(rst), // Global rst DONE
    .clk(clk),// Global clk DONE
    .Register_Destination(Register_Destination), // ptr to register destination from decoder DONE
    .Register_1_operand(Register_1_operand), // ptr to reg1 coming from decoder DONE
    .Register_2_operand(Register_2_operand), // ptr to reg2 coming from decoder DONE
    .RegWrite(RegWrite), // RegWrite comes from FSM DONE
    .data_in(data_in_REG), // Only 2 things that can write to Register file is ALU or RAM load word instruction
    .instr_data_out1(register_1_data), // Outputting reg1 data DONE
    .instr_data_out2(register_2_data) // Outputting reg2 data DONE
    );
    
   
    (* keep_hierarchy = "yes" *)
    RAM Data(
    .clk(clk), // Global Clock DONE
    .write_enable(MemWrite), // Write Enable coming in from FSM DONE
    .address(ALU_Out_Sequential), // Address will come from ALU because the address will be base register 8b address + immediate value for sb and lb DONE
    .data_in(register_1_data), // Register in instruction being stored for sb instructions DONE
    .data_out(RAM_data_out) // RAM data out DONE
    );
    
    assign B = Is_immediate ? extended_immediate : register_2_data; // Decides if B should be immediate or register value
    
    assign A = (instr_Opcode == lw || instr_Opcode == sw) ? register_2_data : register_1_data; // Decides if  A is register 2 data or register 1 data
    
    (* keep_hierarchy = "yes" *)
    ALU Arithmitic(
    .clk(clk),
    .rst(rst),
    .A(A),// source will be driven by lw, sw, or register 1 data DONE
    .B(B), // will be driven by extended signed, unsigned immediate, register value, DONE
    .ALU_Enable(ALU_Enable),
    .ALU_OP(ALUOp), // Taking in ALU_OP from FSM DONE
    .ALU_Out_Sequential(ALU_Out_Sequential), // going out to register file DONE
    .overflow(overflow), // tells us if overflow has occurred, value is valid or not. DONE
    .less_than_flag(less_than_flag), // outputting less than flag DONE
    .is_equal(is_equal), // outputting equal flag DONE
    .zero_flag(zero_flag), // outputting zero flag DONE
    .HI(HI), // upper bits of multiplication instruction DONE
    .LO(LO) // lower bits of multipllication instruction DONE
    );
   
    
    //Top level assignments for simulation
    
    // Top Level FETCH
    assign Current_fetch = Fetch;
    
    // Probing instruction register content in top level module
    assign REG1 = register_1_data;
    assign REG2 = register_2_data;
    
    // Probing FSM state register in top level
    assign Current_state = State; 
    assign IRWrite_Top = IRWrite;
    assign MemWrite_Top = MemWrite;
    assign MemRead_Top = MemRead;
    assign PC_en_Top = PC_en;
    assign RegWrite_Top = RegWrite;
    
    // Probing PC in top level
    assign PC = pc;
    
    // Probing ALU_out for top level module
    assign ALU_Data = ALU_Out_Sequential; 
    
  
 //FOR TESTBENCHING SIMULATION ONLY  
reg [80*8:1] opcode_name;  // string

always @(*) begin
    case (instr_Opcode)
        addi: opcode_name = "ADDI";
        add : opcode_name = "ADD";
        lw  : opcode_name = "LW";
        subi: opcode_name = "SUBI";
        sub : opcode_name = "SUB";
        beq : opcode_name = "BEQ";
        bne : opcode_name = "BNE";
        slt : opcode_name = "SLT";
        slti: opcode_name = "SLTI";
        jump: opcode_name = "JUMP";
        sw  : opcode_name = "SW";
        sra : opcode_name = "SRA";
        sll : opcode_name = "SLL";
        HLT : opcode_name = "HLT";
        default: opcode_name = "UNKNOWN";
    endcase
end

always @(posedge clk) begin
    $display("T=%0t | PC=%0d | Fetch=%h | State=%0d | Instruction =%0s | ALUsrcA = %0d | ALUsrcB = %0d |ALU_Out = %0d | IRwrite = %0d | Regwrite = %0d | Register Destination = %0d | Instruction Register 1 data = %0d | Instruction Register 2 data = %0d",
             $time, pc, Fetch, State, opcode_name,A,B,ALU_Out_Sequential,IRWrite,RegWrite,Register_Destination,register_1_data,register_2_data);
end




endmodule
